----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity FIFO is
	port (
			clk :in  std_logic;
			dataout  : out std_logic_vector (7 downto 0);
			dataout2 : out std_logic_vector (7 downto 0);
			led: out std_logic_vector(3 downto 0);
			Rx: in std_logic;
			Tx: out std_logic
			);
end FIFO;

architecture Behavioral of FIFO is
	
TYPE State_type IS (empezar,empezar11,empezar21,empezar31,empezar41, apagar, reiniciar, salir,fempezar,
fempezar11,fempezar21,fempezar31,fempezar41, fapagar, freiniciar, fsalir, espera); 
SIGNAL State : State_Type; 
signal contador: integer range 0 to 12800;
signal flag: std_logic;
signal contbit: integer range 0 to 1250;
signal num: integer range 0 to 10;
signal vector: std_logic_vector (7 downto 0);
signal enable11: std_logic:='0';
signal enable21: std_logic:='0';
signal enable31: std_logic:='0';
signal enable41: std_logic:='0';
signal bits: integer range 0 to 15:=0;
signal tiempo: integer range 0 to 11999999:=0;
	
	signal i,i1,i2,i3 : integer range 0 to 99:=0;
	
		type memory_type is array (0 to 99) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
	signal sine : memory_type :=(  254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 2, 1, 0, 0, 0, 1, 2, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253);
		signal trian : memory_type :=(255, 250, 245, 240, 235, 230,
											  	225, 220, 215, 210, 205, 200,
											  	195, 190, 185, 180, 175, 170,
										     	165, 160, 155, 150, 145, 140, 
											  	135, 130, 125, 120, 115, 110, 
											 	100, 95,  90, 85, 80, 75, 70,
											  	65, 60, 55, 50, 45, 40, 35, 30,
											  	25, 20, 15, 10, 5, 0, 0, 5,
											  	10, 15, 20, 25, 30, 35, 40,
											  	45, 50, 55, 60, 65, 70, 75, 80,
											  	85, 90, 95, 100, 105, 110, 115, 
											  	120, 125, 130, 135, 140, 145, 150, 
											  	155, 160, 165, 170, 175, 180,
											  	185, 190, 195, 200, 205, 210,
											  	215, 220, 225, 230, 235, 240);
	signal triansie : memory_type :=(255, 0, 5, 10, 15, 20,
												25, 30, 35, 40, 45, 50, 55, 60,
												65, 70, 75, 80,85, 90, 95, 100,
												105, 110, 115, 120, 125, 130,
												135, 145, 150, 155, 160, 165,
												170, 175, 180, 185, 190, 200,
												250, 0, 5, 10, 15, 20, 25,
												30, 35, 40, 45, 50, 55, 60, 65,
												70, 75, 80, 85, 90, 95, 100, 105,
												110, 115, 120, 125, 130, 135, 140, 145,
												150, 155, 160, 165, 170, 175, 180, 185,
												190, 195, 200, 205, 230, 235, 240, 245, 
												250, 255, 0, 5, 10, 15, 20, 25, 30, 35,
												40, 45, 50);
	signal gauss : memory_type :=(  0,0,0, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253, 254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 0, 0, 0,0);
			
begin
process(clk)
begin
--to check the rising edge of the clock signal
if(rising_edge(clk)) then 
if rx = '0' then
		flag <= '1';
	end if;
	if flag = '1' then
		if contador = 12800 then 
			contador <= 0;
			flag <= '0';
			num <= 0;
		elsif contador = 0 and rx = '0' then
			contador <= contador + 1;
		else 
			contador <= contador + 1;
			if contbit = 1249 then
				num <= num + 1;
				contbit <= 0;
			else contbit <= contbit + 1;
			end if;
		end if;
	end if;
	
	Case num is
		when 1 => vector(0) <= rx;
		when 2 => vector(1) <= rx;
		when 3 => vector(2) <= rx;
		when 4 => vector(3) <= rx;
		when 5 => vector(4) <= rx;
		when 6 => vector(5) <= rx;
		when 7 => vector(6) <= rx;
      when 8 => vector(7) <= rx;		
		when others => tx<= rx ;
	end case;
	
	tx <= rx;

case state is 

	when espera =>
		case vector is
			when "00110001" => ----1
				state<=empezar;
			when "00110010" => ----2
				state<=apagar;
			when "00110011" => ----3
				state<=reiniciar;
			when "00110100" => ----4
				state<=salir;
			when "00110101" => ----5
				state<=empezar11;
			when "00110110" => ----6
				state<=empezar21;
			when "00110111" => ----7
				state<=empezar31;
			when "00111000" => ----8
				state<=empezar41;
			when others =>
				state<=espera;
		end case;
		
	when empezar11 =>
		enable11 <= '1';
		enable21 <= '0';
		enable31 <= '0';
		enable41 <= '0';
		state <= fempezar11;
	when fempezar11 =>
		if vector /= "00110101" then
			state<=espera;
		else 
			state<=fempezar11;
		end if;
		
	when empezar21 =>
		enable11 <= '0';
		enable21 <= '1';
		enable31 <= '0';
		enable41 <= '0';
		state <= fempezar21;
	when fempezar21 =>
		if vector /= "00110110" then
			state<=espera;
		else 
			state<=fempezar21;
		end if;
		
	when empezar31 =>
		enable11 <= '0';
		enable21 <= '0';
		enable31 <= '1';
		enable41 <= '0';
		state <= fempezar31;
	when fempezar31 =>
		if vector /= "00110111" then
			state<=espera;
		else 
			state<=fempezar31;
		end if;

	when empezar41 =>
		enable11 <= '0';
		enable21 <= '0';
		enable31 <= '0';
		enable41 <= '1';
		state <= fempezar41;
	when fempezar41 =>
		if vector /= "00111000" then
			state<=espera;
		else 
			state<=fempezar41;
		end if;
		
	when apagar =>
		enable11 <= '0';
		enable21 <= '0';
		enable31 <= '0';
		enable41 <= '0';
		state <=fapagar;
	when fapagar =>
		if vector /= "00110010" then
			state<=espera;
		else 
			state<=fapagar;
		end if;
		
	when reiniciar =>
		i<=0;
		i1<=0;
		i2<=0;
		i3<=0;
		tiempo<=0;
		state <=freiniciar;
	when freiniciar =>
		if vector /= "00110011" then
			state<=espera;
		else 
			state<=freiniciar;
		end if;	
		
	when salir =>
		enable11<='0';
		enable21<='0';
		enable31<='0';
		enable41<='0';
		i<=0;
		i1<=0;
		i2<=0;
		i3<=0;
		dataout <= std_logic_vector(to_unsigned(sine(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sine(0),8));
		dataout2 <= std_logic_vector(to_unsigned(trian(0),8));
		dataout2 <= std_logic_vector(to_unsigned(triansie(0),8));
		dataout2 <= std_logic_vector(to_unsigned(gauss(0),8));
		state <=fsalir;
	when fsalir =>
		if vector /= "00110100" then
			state<=espera;
		else 
			state<=fsalir;
		end if;	
		
	when others =>
		state<=espera;	
end case;	
	
	if enable11 = '1' then
		dataout <= std_logic_vector(to_unsigned(sine(i),8));
		dataout2 <= std_logic_vector(to_unsigned(sine(i),8));
		i <= i+ 1;
			if(i = 99) then
			i <= 0;
			end if;
	end if;
	
	if enable21 = '1' then
		dataout2 <= std_logic_vector(to_unsigned((trian(i1)),8));
		i1 <= i1 + 1;
		if(i1 = 99) then
			i1 <= 0;
		end if;
	end if;

	if enable31 = '1' then
		dataout2 <= std_logic_vector(to_unsigned((triansie(i2)),8));
		i2 <= i2 + 1;
		if(i2 = 99) then
			i2 <= 0;
		end if;
	end if;
	
		if enable41 = '1' then
		dataout2 <= std_logic_vector(to_unsigned((gauss(i3)),8));
		i3 <= i3 + 1;
	end if;
				
end if;
end process;					
end Behavioral;
