----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity FIFO is
	port (
			clk :in  std_logic;
			dataout  : out std_logic_vector (7 downto 0);
			dataout2 : out std_logic_vector (7 downto 0);
			led: out std_logic_vector(3 downto 0);
			Rx: in std_logic;
			Tx: out std_logic
			);
end FIFO;

architecture Behavioral of FIFO is
	
TYPE State_type IS (apagar, reiniciar, salir,fapagar, freiniciar, fsalir, espera,
empezar111,empezar211,empezar311,empezar411,fempezar111,fempezar211,fempezar311,fempezar411,
empezar112,empezar212,empezar312,empezar412,fempezar112,fempezar212,fempezar312,fempezar412,
empezar113,empezar213,empezar313,empezar413,fempezar113,fempezar213,fempezar313,fempezar413,
empezar121,empezar221,empezar321,empezar421,fempezar121,fempezar221,fempezar321,fempezar421,
empezar122,empezar222,empezar322,empezar422,fempezar122,fempezar222,fempezar322,fempezar422,
empezar123,empezar223,empezar323,empezar423,fempezar123,fempezar223,fempezar323,fempezar423);

SIGNAL State : State_Type; 
signal contador: integer range 0 to 12800;
signal flag: std_logic;
signal contbit: integer range 0 to 1250;
signal num: integer range 0 to 10;
signal vector: std_logic_vector (7 downto 0);

signal enable111: std_logic:='0';
signal enable211: std_logic:='0';
signal enable311: std_logic:='0';
signal enable411: std_logic:='0';

signal enable112: std_logic:='0';
signal enable212: std_logic:='0';
signal enable312: std_logic:='0';
signal enable412: std_logic:='0';

signal enable113: std_logic:='0';
signal enable213: std_logic:='0';
signal enable313: std_logic:='0';
signal enable413: std_logic:='0';

signal enable121: std_logic:='0';
signal enable221: std_logic:='0';
signal enable321: std_logic:='0';
signal enable421: std_logic:='0';

signal enable122: std_logic:='0';
signal enable222: std_logic:='0';
signal enable322: std_logic:='0';
signal enable422: std_logic:='0';

signal enable123: std_logic:='0';
signal enable223: std_logic:='0';
signal enable323: std_logic:='0';
signal enable423: std_logic:='0';

signal bits: integer range 0 to 15:=0;
signal tiempo: integer range 0 to 11999999:=0;

	signal i,i1,i2,i3 : integer range 0 to 99:=0;
	signal j,j1,j2,j3 : integer range 0 to 99:=0;
	signal k,k1,k2,k3 : integer range 0 to 99:=0;
	signal l,l1,l2,l3 : integer range 0 to 99:=0;
	signal m,m1,m2,m3 : integer range 0 to 99:=0;
	signal n,n1,n2,n3 : integer range 0 to 99:=0;
	
		type memory_type is array (0 to 99) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
	signal sine11 : memory_type :=(254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 2, 1, 0, 0, 0, 1, 2, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253);
		signal trian11 : memory_type :=(255, 250, 245, 240, 235, 230,
											  	225, 220, 215, 210, 205, 200,
											  	195, 190, 185, 180, 175, 170,
										     	165, 160, 155, 150, 145, 140, 
											  	135, 130, 125, 120, 115, 110, 
											 	100, 95,  90, 85, 80, 75, 70,
											  	65, 60, 55, 50, 45, 40, 35, 30,
											  	25, 20, 15, 10, 5, 0, 0, 5,
											  	10, 15, 20, 25, 30, 35, 40,
											  	45, 50, 55, 60, 65, 70, 75, 80,
											  	85, 90, 95, 100, 105, 110, 115, 
											  	120, 125, 130, 135, 140, 145, 150, 
											  	155, 160, 165, 170, 175, 180,
											  	185, 190, 195, 200, 205, 210,
											  	215, 220, 225, 230, 235, 240);
	signal sierra11 : memory_type :=(255, 0, 5, 10, 15, 20,
												25, 30, 35, 40, 45, 50, 55, 60,
												65, 70, 75, 80,85, 90, 95, 100,
												105, 110, 115, 120, 125, 130,
												135, 145, 150, 155, 160, 165,
												170, 175, 180, 185, 190, 200,
												250, 0, 5, 10, 15, 20, 25,
												30, 35, 40, 45, 50, 55, 60, 65,
												70, 75, 80, 85, 90, 95, 100, 105,
												110, 115, 120, 125, 130, 135, 140, 145,
												150, 155, 160, 165, 170, 175, 180, 185,
												190, 195, 200, 205, 230, 235, 240, 245, 
												250, 255, 0, 5, 10, 15, 20, 25, 30, 35,
												40, 45, 50);
	signal gauss11 : memory_type :=(0,0,0, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253, 254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 0, 0, 0,0);
		type memory_type2 is array (0 to 99) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
	signal sine12 : memory_type2 :=(50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8, 10, 15, 19, 24, 27, 34, 42,
												50, 50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8, 10, 15, 19, 24, 27, 34, 42,
												50, 50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8, 10, 15, 19, 24, 27, 34, 42,
												50,50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8);
	signal trian12 : memory_type2 :=(150, 140, 130, 120,
												110, 100, 90, 80, 70, 60, 50, 40, 
												30, 20, 10, 0, 10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150, 140,
												130, 120, 110, 100, 90, 80, 70,
												60, 50, 40, 30, 20, 10, 0, 10,
												20, 30, 40, 50, 60, 70, 80, 90, 100,
												110, 120, 130, 140, 150, 140, 130, 120,
												110, 100, 90, 80, 70, 60, 50, 40, 
												30, 20, 10, 0,
												10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150, 140,
												130, 120, 110, 100, 90, 80, 70, 60);
	signal sierra12 : memory_type2 :=(0, 10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150,
												0, 10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150,
												0, 10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150,
												0, 10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150,
												0, 10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150,
												0, 10, 20, 30, 40, 50, 60, 70, 80,
												90, 100, 110, 120, 130, 140, 150,
												0, 10, 20, 30);
	signal gauss12 : memory_type2 :=(0,0,0, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253, 254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 0, 0, 0,0);
		type memory_type3 is array (0 to 99) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
	signal sine13 : memory_type3 :=(50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8, 10, 15, 19, 24, 27, 34, 42,
												50, 50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8, 10, 15, 19, 24, 27, 34, 42,
												50, 50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8, 10, 15, 19, 24, 27, 34, 42,
												50,50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8);
	signal trian13 : memory_type3 :=(255, 250, 245, 240, 235, 230,
											  	225, 220, 215, 210, 205, 200,
											  	195, 190, 185, 180, 175, 170,
										     	165, 160, 155, 150, 145, 140, 
											  	135, 130, 125, 120, 115, 110, 
											 	100, 95,  90, 85, 80, 75, 70,
											  	65, 60, 55, 50, 45, 40, 35, 30,
											  	25, 20, 15, 10, 5, 0, 0, 5,
											  	10, 15, 20, 25, 30, 35, 40,
											  	45, 50, 55, 60, 65, 70, 75, 80,
											  	85, 90, 95, 100, 105, 110, 115, 
											  	120, 125, 130, 135, 140, 145, 150, 
											  	155, 160, 165, 170, 175, 180,
											  	185, 190, 195, 200, 205, 210,
											  	215, 220, 225, 230, 235, 240);
	signal sierra13 : memory_type3 :=(255, 0, 5, 10, 15, 20,
												25, 30, 35, 40, 45, 50, 55, 60,
												65, 70, 75, 80,85, 90, 95, 100,
												105, 110, 115, 120, 125, 130,
												135, 145, 150, 155, 160, 165,
												170, 175, 180, 185, 190, 200,
												250, 0, 5, 10, 15, 20, 25,
												30, 35, 40, 45, 50, 55, 60, 65,
												70, 75, 80, 85, 90, 95, 100, 105,
												110, 115, 120, 125, 130, 135, 140, 145,
												150, 155, 160, 165, 170, 175, 180, 185,
												190, 195, 200, 205, 230, 235, 240, 245, 
												250, 255, 0, 5, 10, 15, 20, 25, 30, 35,
												40, 45, 50);
	signal gauss13 : memory_type3 :=(0,0,0, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253, 254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 0, 0, 0,0);
		type memory_type4 is array (0 to 99) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
	signal sine21 : memory_type4 :=(27, 34, 42, 50, 58, 66, 
												73, 81, 88, 95, 101, 107,												
												113, 119, 124, 129, 134, 138,
												141, 145, 147, 150, 150,
												147, 145, 141, 138, 134, 129,
												124, 119, 113, 107, 101, 95, 88, 81, 
												73, 66, 58, 50, 42, 34, 27, 24, 
												19, 15, 10, 8, 6, 3, 1, 0, 0, 1, 2, 3, 6,
												8, 10, 15, 19, 24, 27, 34, 42,
												50, 58, 66, 73, 81, 88, 195,
												101, 101, 107, 113, 119, 124, 129, 134, 138,
												141, 145, 147, 150, 150,
												147, 145, 141, 138, 134, 129,
												124, 119, 113, 107, 101, 95, 88);
	signal trian21 : memory_type4 :=(255, 250, 245, 240, 235, 230,
											  	225, 220, 215, 210, 205, 200,
											  	195, 190, 185, 180, 175, 170,
										     	165, 160, 155, 150, 145, 140, 
											  	135, 130, 125, 120, 115, 110, 
											 	100, 95,  90, 85, 80, 75, 70,
											  	65, 60, 55, 50, 45, 40, 35, 30,
											  	25, 20, 15, 10, 5, 0, 0, 5,
											  	10, 15, 20, 25, 30, 35, 40,
											  	45, 50, 55, 60, 65, 70, 75, 80,
											  	85, 90, 95, 100, 105, 110, 115, 
											  	120, 125, 130, 135, 140, 145, 150, 
											  	155, 160, 165, 170, 175, 180,
											  	185, 190, 195, 200, 205, 210,
											  	215, 220, 225, 230, 235, 240);
	signal sierra21 : memory_type4 :=(255, 0, 5, 10, 15, 20,
												25, 30, 35, 40, 45, 50, 55, 60,
												65, 70, 75, 80,85, 90, 95, 100,
												105, 110, 115, 120, 125, 130,
												135, 145, 150, 155, 160, 165,
												170, 175, 180, 185, 190, 200,
												250, 0, 5, 10, 15, 20, 25,
												30, 35, 40, 45, 50, 55, 60, 65,
												70, 75, 80, 85, 90, 95, 100, 105,
												110, 115, 120, 125, 130, 135, 140, 145,
												150, 155, 160, 165, 170, 175, 180, 185,
												190, 195, 200, 205, 230, 235, 240, 245, 
												250, 255, 0, 5, 10, 15, 20, 25, 30, 35,
												40, 45, 50);
	signal gauss21 : memory_type4 :=(0,0,0, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253, 254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 0, 0, 0,0);
		type memory_type5 is array (0 to 99) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
	signal sine22 : memory_type5 :=(254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 2, 1, 0, 0, 0, 1, 2, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253);
	signal trian22 : memory_type5 :=(255, 250, 245, 240, 235, 230,
											  	225, 220, 215, 210, 205, 200,
											  	195, 190, 185, 180, 175, 170,
										     	165, 160, 155, 150, 145, 140, 
											  	135, 130, 125, 120, 115, 110, 
											 	100, 95,  90, 85, 80, 75, 70,
											  	65, 60, 55, 50, 45, 40, 35, 30,
											  	25, 20, 15, 10, 5, 0, 0, 5,
											  	10, 15, 20, 25, 30, 35, 40,
											  	45, 50, 55, 60, 65, 70, 75, 80,
											  	85, 90, 95, 100, 105, 110, 115, 
											  	120, 125, 130, 135, 140, 145, 150, 
											  	155, 160, 165, 170, 175, 180,
											  	185, 190, 195, 200, 205, 210,
											  	215, 220, 225, 230, 235, 240);
	signal sierra22 : memory_type5 :=(255, 0, 5, 10, 15, 20,
												25, 30, 35, 40, 45, 50, 55, 60,
												65, 70, 75, 80,85, 90, 95, 100,
												105, 110, 115, 120, 125, 130,
												135, 145, 150, 155, 160, 165,
												170, 175, 180, 185, 190, 200,
												250, 0, 5, 10, 15, 20, 25,
												30, 35, 40, 45, 50, 55, 60, 65,
												70, 75, 80, 85, 90, 95, 100, 105,
												110, 115, 120, 125, 130, 135, 140, 145,
												150, 155, 160, 165, 170, 175, 180, 185,
												190, 195, 200, 205, 230, 235, 240, 245, 
												250, 255, 0, 5, 10, 15, 20, 25, 30, 35,
												40, 45, 50);
	signal gauss22 : memory_type5 :=(0,0,0, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253, 254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 0, 0, 0,0);
		type memory_type6 is array (0 to 99) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
	signal sine23 : memory_type6 :=(254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 2, 1, 0, 0, 0, 1, 2, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253);
	signal trian23 : memory_type6 :=(255, 250, 245, 240, 235, 230,
											  	225, 220, 215, 210, 205, 200,
											  	195, 190, 185, 180, 175, 170,
										     	165, 160, 155, 150, 145, 140, 
											  	135, 130, 125, 120, 115, 110, 
											 	100, 95,  90, 85, 80, 75, 70,
											  	65, 60, 55, 50, 45, 40, 35, 30,
											  	25, 20, 15, 10, 5, 0, 0, 5,
											  	10, 15, 20, 25, 30, 35, 40,
											  	45, 50, 55, 60, 65, 70, 75, 80,
											  	85, 90, 95, 100, 105, 110, 115, 
											  	120, 125, 130, 135, 140, 145, 150, 
											  	155, 160, 165, 170, 175, 180,
											  	185, 190, 195, 200, 205, 210,
											  	215, 220, 225, 230, 235, 240);
	signal sierra23 : memory_type6 :=(255, 0, 5, 10, 15, 20,
												25, 30, 35, 40, 45, 50, 55, 60,
												65, 70, 75, 80,85, 90, 95, 100,
												105, 110, 115, 120, 125, 130,
												135, 145, 150, 155, 160, 165,
												170, 175, 180, 185, 190, 200,
												250, 0, 5, 10, 15, 20, 25,
												30, 35, 40, 45, 50, 55, 60, 65,
												70, 75, 80, 85, 90, 95, 100, 105,
												110, 115, 120, 125, 130, 135, 140, 145,
												150, 155, 160, 165, 170, 175, 180, 185,
												190, 195, 200, 205, 230, 235, 240, 245, 
												250, 255, 0, 5, 10, 15, 20, 25, 30, 35,
												40, 45, 50);
	signal gauss23 : memory_type6 :=(0,0,0, 3, 6,
												8, 12, 15, 19, 24, 29, 34, 40,
												46, 52, 58, 65, 72, 80, 87, 95,
												103, 111, 119, 127, 134, 142, 150, 158, 166, 
												173, 181, 188, 195, 201, 207,
												213, 219, 224, 229, 234, 238,
												241, 245, 247, 250, 251, 252, 
												253, 254, 253, 252, 251, 250,
											  247, 245, 241, 238, 234, 229,
											  224, 219, 213, 207, 201, 195,
												188, 181, 173, 166, 158, 150,
												142, 134, 127, 119, 111, 103,
												95, 87, 80, 72, 65, 58, 52, 46, 
												40, 34, 29, 24, 19, 15, 12, 8, 
												6, 3, 0, 0, 0,0);
			
begin
process(clk)
begin
--to check the rising edge of the clock signal
if(rising_edge(clk)) then 
if rx = '0' then
		flag <= '1';
	end if;
	if flag = '1' then
		if contador = 12800 then 
			contador <= 0;
			flag <= '0';
			num <= 0;
		elsif contador = 0 and rx = '0' then
			contador <= contador + 1;
		else 
			contador <= contador + 1;
			if contbit = 1249 then
				num <= num + 1;
				contbit <= 0;
			else contbit <= contbit + 1;
			end if;
		end if;
	end if;
	
	Case num is
		when 1 => vector(0) <= rx;
		when 2 => vector(1) <= rx;
		when 3 => vector(2) <= rx;
		when 4 => vector(3) <= rx;
		when 5 => vector(4) <= rx;
		when 6 => vector(5) <= rx;
		when 7 => vector(6) <= rx;
      when 8 => vector(7) <= rx;		
		when others => tx<= rx ;
	end case;
	
	tx <= rx;

case state is 

	when espera =>
		case vector is
			when "00110000" => ----0
				state<=salir;
			when "00110001" => ----1
				state<=reiniciar;
			when "00110010" => ----2
				state<=empezar111;
			when "00110011" => ----3
				state<=empezar211;
			when "00110100" => ----4
				state<=empezar311;
			when "00110101" => ----5
				state<=empezar411;
			when "00110110" => ----6
				state<=empezar112;
			when "00110111" => ----7
				state<=empezar212;
			when "00111000" => ----8
				state<=empezar312;
			when "00111001" => ----9
				state<=empezar412;
			when "00111010" => ----10
				state<=empezar113;
			when "00111011" => ----11
				state<=empezar213;
			when "00111100" => ----12
				state<=empezar313;
			when "00111101" => ----13
				state<=empezar413;
			when "00111110" => ----14
				state<=empezar121;
			when "00111111" => ----15
				state<=empezar221;
			when others =>
				state<=salir;
		end case;
		
	when salir =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		i<=0;
		i1<=0;
		i2<=0;
		i3<=0;
		j<=0;
		j1<=0;
		j2<=0;
		j3<=0;
		k<=0;
		k1<=0;
		k2<=0;
		k3<=0;
		m<=0;		
		l<=0;
		l1<=0;
		l2<=0;
		l3<=0;
		m<=0;
		m1<=0;
		m2<=0;
		m3<=0;
		n<=0;
		n1<=0;
		n2<=0;
		n3<=0;
		dataout2 <= std_logic_vector(to_unsigned(sine11(0),8));
		dataout2 <= std_logic_vector(to_unsigned(trian11(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sierra11(0),8));
		dataout2 <= std_logic_vector(to_unsigned(gauss11(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sine12(0),8));
		dataout2 <= std_logic_vector(to_unsigned(trian12(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sierra12(0),8));
		dataout2 <= std_logic_vector(to_unsigned(gauss12(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sine13(0),8));
		dataout2 <= std_logic_vector(to_unsigned(trian13(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sierra13(0),8));
		dataout2 <= std_logic_vector(to_unsigned(gauss13(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sine21(0),8));
		dataout2 <= std_logic_vector(to_unsigned(trian21(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sierra21(0),8));
		dataout2 <= std_logic_vector(to_unsigned(gauss21(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sine22(0),8));
		dataout2 <= std_logic_vector(to_unsigned(trian22(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sierra22(0),8));
		dataout2 <= std_logic_vector(to_unsigned(gauss22(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sine23(0),8));
		dataout2 <= std_logic_vector(to_unsigned(trian23(0),8));
		dataout2 <= std_logic_vector(to_unsigned(sierra23(0),8));
		dataout2 <= std_logic_vector(to_unsigned(gauss23(0),8));

		state <=fsalir;
	when fsalir =>
		if vector /= "00110000" then
			state<=espera;
		else 
			state<=fsalir;
		end if;

	when reiniciar =>
		i<=0;
		i1<=0;
		i2<=0;
		i3<=0;
		j<=0;
		j1<=0;
		j2<=0;
		j3<=0;
		k<=0;
		k1<=0;
		k2<=0;
		k3<=0;
		l<=0;
		l1<=0;
		l2<=0;
		l3<=0;
		m<=0;
		m1<=0;
		m2<=0;
		m3<=0;
		n<=0;
		n1<=0;
		n2<=0;
		n3<=0;
		tiempo<=0;
		state <=freiniciar;
	when freiniciar =>
		if vector /= "00110001" then
			state<=espera;
		else 
			state<=freiniciar;
		end if;		
	
	when empezar111 =>
		enable111 <= '1';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar111;
	when fempezar111 =>
		if vector /= "00110010" then
			state<=espera;
		else 
			state<=fempezar111;
		end if;
		
	when empezar211 =>
		enable111 <= '0';
		enable211 <= '1';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';		
		state <= fempezar211;
	when fempezar211 =>
		if vector /= "00110011" then
			state<=espera;
		else 
			state<=fempezar211;
		end if;
		
	when empezar311 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '1';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar311;
	when fempezar311 =>
		if vector /= "00110100" then
			state<=espera;
		else 
			state<=fempezar311;
		end if;

	when empezar411 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '1';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar411;
	when fempezar411 =>
		if vector /= "00110101" then
			state<=espera;
		else 
			state<=fempezar411;
		end if;

	when empezar112 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '1';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar112;
	when fempezar112 =>
		if vector /= "00110110" then
			state<=espera;
		else 
			state<=fempezar112;
		end if;
		
	when empezar212 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '1';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';		
		state <= fempezar212;
	when fempezar212 =>
		if vector /= "00110111" then
			state<=espera;
		else 
			state<=fempezar212;
		end if;
		
	when empezar312 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '1';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar312;
	when fempezar312 =>
		if vector /= "00111000" then
			state<=espera;
		else 
			state<=fempezar312;
		end if;

	when empezar412 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '1';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar412;
	when fempezar412 =>
		if vector /= "00111001" then
			state<=espera;
		else 
			state<=fempezar412;
		end if;
		
	when empezar113 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '1';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar113;
	when fempezar113 =>
		if vector /= "00111010" then
			state<=espera;
		else 
			state<=fempezar113;
		end if;
		
	when empezar213 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '1';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';		
		state <= fempezar213;
	when fempezar213 =>
		if vector /= "00111011" then
			state<=espera;
		else 
			state<=fempezar213;
		end if;
		
	when empezar313 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '1';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar313;
	when fempezar313 =>
		if vector /= "00111100" then
			state<=espera;
		else 
			state<=fempezar313;
		end if;

	when empezar413 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '1';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar413;
	when fempezar413 =>
		if vector /= "00111101" then
			state<=espera;
		else 
			state<=fempezar413;
		end if;

	when empezar121 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '1';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar121;
	when fempezar121 =>
		if vector /= "00111110" then
			state<=espera;
		else 
			state<=fempezar121;
		end if;
		
	when empezar221 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '1';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';		
		state <= fempezar221;
	when fempezar221 =>
		if vector /= "00111111" then
			state<=espera;
		else 
			state<=fempezar221;
		end if;
		
	when empezar321 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '1';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar321;
	when fempezar321 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar321;
		end if;

	when empezar421 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '1';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar421;
	when fempezar421 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar421;
		end if;

	when empezar122 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '1';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar122;
	when fempezar122 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar122;
		end if;
		
	when empezar222 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '1';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';		
		state <= fempezar222;
	when fempezar222 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar222;
		end if;
		
	when empezar322 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '1';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar322;
	when fempezar322 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar322;
		end if;

	when empezar422 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '1';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar422;
	when fempezar422 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar422;
		end if;

	when empezar123 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '1';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '0';
		state <= fempezar123;
	when fempezar123 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar123;
		end if;
		
	when empezar223 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '1';
		enable323 <= '0';
		enable423 <= '0';		
		state <= fempezar223;
	when fempezar223 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar223;
		end if;
		
	when empezar323 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '1';
		enable423 <= '0';
		state <= fempezar323;
	when fempezar323 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar323;
		end if;

	when empezar423 =>
		enable111 <= '0';
		enable211 <= '0';
		enable311 <= '0';
		enable411 <= '0';
		enable112 <= '0';
		enable212 <= '0';
		enable312 <= '0';
		enable412 <= '0';
		enable113 <= '0';
		enable213 <= '0';
		enable313 <= '0';
		enable413 <= '0';
		enable121 <= '0';
		enable221 <= '0';
		enable321 <= '0';
		enable421 <= '0';
		enable122 <= '0';
		enable222 <= '0';
		enable322 <= '0';
		enable422 <= '0';
		enable123 <= '0';
		enable223 <= '0';
		enable323 <= '0';
		enable423 <= '1';
		state <= fempezar423;
	when fempezar423 =>
		if vector /= "" then
			state<=espera;
		else 
			state<=fempezar423;
		end if;
		
	when others =>
		state<=espera;	
end case;	
	
	if enable111 = '1' then
		dataout <= std_logic_vector(to_unsigned(sine11(i),8));
		dataout2 <= std_logic_vector(to_unsigned(sine11(i),8));
		i <= i+ 1;
			if(i = 99) then
			i <= 0;
			end if;
	end if;
	
	if enable211 = '1' then
		dataout <= std_logic_vector(to_unsigned(trian11(i1),8));
		dataout2 <= std_logic_vector(to_unsigned((trian11(i1)),8));
		i1 <= i1 + 1;
		if(i1 = 99) then
			i1 <= 0;
		end if;
	end if;

	if enable311 = '1' then
		dataout <= std_logic_vector(to_unsigned(sierra11(i2),8));
		dataout2 <= std_logic_vector(to_unsigned((sierra11(i2)),8));
		i2 <= i2 + 1;
		if(i2 = 99) then
			i2 <= 0;
		end if;
	end if;
	
		if enable411 = '1' then
		dataout <= std_logic_vector(to_unsigned(gauss11(i3),8));
		dataout2 <= std_logic_vector(to_unsigned((gauss11(i3)),8));
		i3 <= i3 + 1;
	end if;
	
	if enable112 = '1' then
		dataout <= std_logic_vector(to_unsigned(sine12(j),8));
		dataout2 <= std_logic_vector(to_unsigned(sine12(j),8));
		j <= j+ 1;
			if(j = 99) then
			j <= 0;
			end if;
	end if;
	
	if enable212 = '1' then
		dataout <= std_logic_vector(to_unsigned(trian12(j1),8));
		dataout2 <= std_logic_vector(to_unsigned((trian12(j1)),8));
		j1 <= j1 + 1;
		if(j1 = 99) then
			j1 <= 0;
		end if;
	end if;

	if enable312 = '1' then
		dataout <= std_logic_vector(to_unsigned(sierra12(j2),8));
		dataout2 <= std_logic_vector(to_unsigned((sierra12(j2)),8));
		j2 <= j2 + 1;
		if(j2 = 99) then
			j2 <= 0;
		end if;
	end if;
	
		if enable412 = '1' then
		dataout <= std_logic_vector(to_unsigned(gauss12(j3),8));
		dataout2 <= std_logic_vector(to_unsigned((gauss12(j3)),8));
		j3 <= j3 + 1;
	end if;
	
	if enable113 = '1' then
		dataout <= std_logic_vector(to_unsigned(sine13(k),8));
		dataout2 <= std_logic_vector(to_unsigned(sine13(k),8));
		k <= k+ 1;
			if(k = 99) then
			k <= 0;
			end if;
	end if;
	
	if enable212 = '1' then
		dataout <= std_logic_vector(to_unsigned(trian13(k1),8));
		dataout2 <= std_logic_vector(to_unsigned((trian13(k1)),8));
		k1 <= k1 + 1;
		if(k1 = 99) then
			k1 <= 0;
		end if;
	end if;

	if enable313 = '1' then
		dataout <= std_logic_vector(to_unsigned(sierra13(k2),8));
		dataout2 <= std_logic_vector(to_unsigned((sierra13(k2)),8));
		k2 <= k2 + 1;
		if(k2 = 99) then
			k2 <= 0;
		end if;
	end if;
	
		if enable413 = '1' then
		dataout <= std_logic_vector(to_unsigned(gauss13(k3),8));
		dataout2 <= std_logic_vector(to_unsigned((gauss13(k3)),8));
		k3 <= k3 + 1;
	end if;

	if enable121 = '1' then
		dataout <= std_logic_vector(to_unsigned(sine21(l),8));
		dataout2 <= std_logic_vector(to_unsigned(sine21(l),8));
		l <= l+ 1;
			if(l = 99) then
			l <= 0;
			end if;
	end if;
	
	if enable221 = '1' then
		dataout <= std_logic_vector(to_unsigned(trian21(l1),8));
		dataout2 <= std_logic_vector(to_unsigned((trian21(l1)),8));
		l1 <= l1 + 1;
		if(l1 = 99) then
			l1 <= 0;
		end if;
	end if;

	if enable321 = '1' then
		dataout <= std_logic_vector(to_unsigned(sierra21(l2),8));
		dataout2 <= std_logic_vector(to_unsigned((sierra21(l2)),8));
		l2 <= l2 + 1;
		if(l2 = 99) then
			l2 <= 0;
		end if;
	end if;
	
		if enable421 = '1' then
		dataout <= std_logic_vector(to_unsigned(gauss21(l3),8));
		dataout2 <= std_logic_vector(to_unsigned((gauss21(l3)),8));
		l3 <= l3 + 1;
	end if;

	if enable122 = '1' then
		dataout <= std_logic_vector(to_unsigned(sine22(m),8));
		dataout2 <= std_logic_vector(to_unsigned(sine22(m),8));
		m <= m+ 1;
			if(m = 99) then
			m <= 0;
			end if;
	end if;
	
	if enable222 = '1' then
		dataout <= std_logic_vector(to_unsigned(trian22(m1),8));
		dataout2 <= std_logic_vector(to_unsigned((trian22(m1)),8));
		m1 <= m1 + 1;
		if(m1 = 99) then
			m1 <= 0;
		end if;
	end if;

	if enable322 = '1' then
		dataout <= std_logic_vector(to_unsigned(sierra22(m2),8));
		dataout2 <= std_logic_vector(to_unsigned((sierra22(m2)),8));
		m2 <= m2 + 1;
		if(m2 = 99) then
			m2 <= 0;
		end if;
	end if;
	
		if enable422 = '1' then
		dataout <= std_logic_vector(to_unsigned(gauss22(m3),8));
		dataout2 <= std_logic_vector(to_unsigned((gauss22(m3)),8));
		m3 <= m3 + 1;
	end if;
	
		if enable123 = '1' then
		dataout <= std_logic_vector(to_unsigned(sine23(n),8));
		dataout2 <= std_logic_vector(to_unsigned(sine23(n),8));
		n <= n+ 1;
			if(n = 99) then
			n <= 0;
			end if;
	end if;
	
	if enable223 = '1' then
		dataout <= std_logic_vector(to_unsigned(trian23(n1),8));
		dataout2 <= std_logic_vector(to_unsigned((trian23(n1)),8));
		n1 <= n1 + 1;
		if(n1 = 99) then
			n1 <= 0;
		end if;
	end if;

	if enable323 = '1' then
		dataout <= std_logic_vector(to_unsigned(sierra23(n2),8));
		dataout2 <= std_logic_vector(to_unsigned((sierra23(n2)),8));
		n2 <= n2 + 1;
		if(n2 = 99) then
			n2 <= 0;
		end if;
	end if;
	
		if enable423 = '1' then
		dataout <= std_logic_vector(to_unsigned(gauss23(n3),8));
		dataout2 <= std_logic_vector(to_unsigned((gauss23(n3)),8));
		n3 <= n3 + 1;
	end if;
	
end if;
end process;					
end Behavioral;